`timescale 1 ns/ 1 ns
module datapath_tb();
reg clk, RST, HALT, MIN_KEY, HR_KEY, INC_SW;
wire[3:0] MS, HOUR;
wire[5:0] SEC, MIN;
wire AMPM;

binary_clock_datapath_rev2 bcdr2(.CLOCK_50(clk),.RST(RST),.HALT(HALT),.MIN_KEY(MIN_KEY),.HR_KEY(HR_KEY),.INC_SW(INC_SW),.ms_out(MS),.sec_out(SEC),.min_out(MIN),.hr_out(HOUR),.AMPM(AMPM));

initial begin
RST <=0; HALT <=0; MIN_KEY <= 1; HR_KEY <= 1; INC_SW <= 0;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
clk <=0; #10; clk <=1; #10;
end
endmodule
 